module tb_spi_fsm;

    

endmodule